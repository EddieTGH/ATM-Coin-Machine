module div_Exception();

endmodule